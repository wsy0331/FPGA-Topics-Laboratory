library IEEE;
use IEEE.std_logic_1164.all;
 
ENTITY pingpong_tb IS
END pingpong_tb;
 
architecture Behavior of pingpong_tb is
    COMPONENT pingpong
        Port (i_clk : in STD_LOGIC;
              i_rst : in STD_LOGIC;
              i_swL : in STD_LOGIC;
              i_swR : in STD_LOGIC;
              o_led : out STD_LOGIC_VECTOR (7 downto 0));
    END COMPONENT;
    
    signal clock : std_logic := '0';
    signal reset : std_logic := '0';
    signal swL : std_logic := '0';
    signal swR : std_logic := '0'; 
    signal led : std_logic_vector(7 downto 0);
    constant clock_period : time := 20 ns;
    
begin
 
    uut: pingpong PORT MAP (
        i_clk => clock,
        i_rst => reset, 
        i_swL => swL,
        i_swR => swR,
        o_led => led
    );    
    
    clock_process :process
    begin
        clock <= '0';
        wait for clock_period/2;
        clock <= '1';
        wait for clock_period/2;
    end process;
    
    stim_proc: process
    begin
        -- ��l�� Reset
        reset <= '0';
        swL <= '0';
        swR <= '0';
        wait for 100 ns;
        reset <= '1';
        wait for 100 ns;
        
        -- Test 1: �k��o�y
        swR <= '1';
        wait for 40 ns;
        swR <= '0';
        wait for 100 ns;
        
        -- Test 2: ���`�若 - ���西�`�^��
        wait for 460 ns;
        swL <= '1';
        wait for 40 ns;
        swL <= '0';
        wait for 100 ns;
        
        -- Test 3: ����S����k��o��
        wait for 460 ns;
        swR <= '1';
        wait for 40 ns;
        swR <= '0';
        wait for 100 ns;
        
        -- Test 4: �k�责�e�� ���b�k���A�B����S����k��o��
        swR <= '1';
        wait for 40 ns;
        swR <= '0';
        wait for 100 ns;
        
        -- Test 5: �k��o�y
        wait for 580 ns;
        swR <= '1';
        wait for 40 ns;
        swR <= '0';
        wait for 100 ns;
        
        -- Test 6: �k��S���쥪��o��
        wait for 860 ns;
        swL <= '1';
        wait for 40 ns;
        swL <= '0';
        wait for 100 ns;   
        
--        --���䴣�e��
--        swL <= '1';
--        wait for 40 ns;
--        swL <= '0';
--        wait for 100 ns;
        
--        --����o�y
--        wait for 460 ns;
--        swL <= '1';
--        wait for 40 ns;
--        swL <= '0';
--        wait for 100 ns;
        
        --�k�䴣����
        wait for 150 ns;
        swR <= '1';
        wait for 40 ns;
        swR <= '0';
        wait for 100 ns;
        
        --����o�y
        wait for 360 ns;
        swL <= '1';
        wait for 40 ns;
        swL <= '0';
        wait for 100 ns;
        
        wait;
    end process;
    
end Behavior;