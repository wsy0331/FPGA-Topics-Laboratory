library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity VGA is
    generic(
        -- 800x600@60Hz SVGA �Ѽ� (40 MHz pixel clock)
        H_RES   : integer   := 800;
        H_FP    : integer   := 40;
        H_SYNC  : integer   := 128;
        H_BP    : integer   := 88;
        H_POL   : std_logic := '1';

        V_RES   : integer   := 600;
        V_FP    : integer   := 1;
        V_SYNC  : integer   := 4;
        V_BP    : integer   := 23;
        V_POL   : std_logic := '1'
    );
    port (
        i_clk    : in  std_logic;  -- 100 MHz System Clock
        i_rst    : in  std_logic;  -- Active-High Reset (Button)
        
        -- Ping Pong Game Inputs
        i_btL    : in  STD_LOGIC;  -- Left Player Button
        i_btR    : in  STD_LOGIC;  -- Right Player Button
        i_swL    : in  STD_LOGIC;  -- Left Player Switch
        i_swR    : in  STD_LOGIC;  -- Right Player Switch
        o_led : out STD_LOGIC_VECTOR (7 downto 0);

        
        -- VGA Outputs
        o_red    : out std_logic_vector(3 downto 0);
        o_green  : out std_logic_vector(3 downto 0);
        o_blue   : out std_logic_vector(3 downto 0);
        o_h_sync : out std_logic;
        o_v_sync : out std_logic
    );
end VGA;

architecture rtl of VGA is

    -- �ޥ� pingpong ����
    component pingpong is
        Port (
            i_clk : in STD_LOGIC;
            i_rst : in STD_LOGIC;  -- active-low
            i_btL : in STD_LOGIC;
            i_btR : in STD_LOGIC;
            i_swL : in STD_LOGIC;
            i_swR : in STD_LOGIC;
            o_led : out STD_LOGIC_VECTOR (7 downto 0)
        );
    end component;

    -- VGA Timing Constants
    constant H_TOTAL : integer := H_RES + H_FP + H_SYNC + H_BP;
    constant V_TOTAL : integer := V_RES + V_FP + V_SYNC + V_BP;

    -- Counters
    signal h_count : integer range 0 to H_TOTAL - 1 := 0;
    signal v_count : integer range 0 to V_TOTAL - 1 := 0;

    -- Pixel Clock Generation (100MHz -> 40MHz)
    signal pix_ce     : std_logic := '0';
    signal ce_idle    : integer range 0 to 3 := 0;
    signal ce_toggle  : std_logic := '0';

    -- Ping Pong Interface Signals
    signal pp_rst_n   : std_logic;              -- Active-low reset for pingpong
    signal led_status : std_logic_vector(7 downto 0); -- Output from pingpong
    
    -- Visual Design Constants (8 "LEDs" on screen)
    constant LED_Y      : integer := 300;       -- Y center position
    constant LED_RADIUS : integer := 30;        -- Radius of the LED circle
    constant LED_GAP    : integer := 90;        -- Horizontal spacing between centers
    constant LED_START_X: integer := 85;        -- X position of the first (left-most) LED
    
begin

    -- Reset Logic: Assuming i_rst is Active-High (1=Reset), 
    -- but pingpong expects Active-Low (0=Reset).
    pp_rst_n <= not i_rst;

    -- ��Ҥ� Ping Pong �C���֤�
    inst_pingpong: pingpong
    port map (
        i_clk => i_clk,
        i_rst => pp_rst_n, -- Convert to active-low
        i_btL => i_btL,
        i_btR => i_btR,
        i_swL => i_swL,
        i_swR => i_swR,
        o_led => led_status
    );

    ------------------------------------------------------------------------
    -- 1. Pixel Clock Enable Generator (100 MHz -> 40 MHz)
    ------------------------------------------------------------------------
    process(i_clk)
    begin
        if rising_edge(i_clk) then
            if i_rst = '1' then
                pix_ce    <= '0';
                ce_idle   <= 0;
                ce_toggle <= '0';
            else
                if ce_idle = 0 then
                    pix_ce <= '1';
                    if ce_toggle = '0' then
                        ce_idle   <= 1;       
                        ce_toggle <= '1';
                    else
                        ce_idle   <= 2;       
                        ce_toggle <= '0';
                    end if;
                else
                    pix_ce  <= '0';
                    ce_idle <= ce_idle - 1;
                end if;
            end if;
        end if;
    end process;

    ------------------------------------------------------------------------
    -- 2. Horizontal Counter
    ------------------------------------------------------------------------
    process(i_clk)
    begin
        if rising_edge(i_clk) then
            if i_rst = '1' then
                h_count <= 0;
            elsif pix_ce = '1' then
                if h_count < H_TOTAL - 1 then
                    h_count <= h_count + 1;
                else
                    h_count <= 0;
                end if;
            end if;
        end if;
    end process;

    ------------------------------------------------------------------------
    -- 3. Vertical Counter
    ------------------------------------------------------------------------
    process(i_clk)
    begin
        if rising_edge(i_clk) then
            if i_rst = '1' then
                v_count <= 0;
            elsif pix_ce = '1' then
                if h_count = H_TOTAL - 1 then
                    if v_count < V_TOTAL - 1 then
                        v_count <= v_count + 1;
                    else
                        v_count <= 0;
                    end if;
                end if;
            end if;
        end if;
    end process;

    ------------------------------------------------------------------------
    -- 4. Sync Signals
    ------------------------------------------------------------------------
    o_h_sync <= H_POL when (h_count >= (H_RES + H_FP) and h_count < (H_RES + H_FP + H_SYNC)) else not H_POL;
    o_v_sync <= V_POL when (v_count >= (V_RES + V_FP) and v_count < (V_RES + V_FP + V_SYNC)) else not V_POL;

    -- 5. RGB Output Logic (Draw 7 Circles based on led_status)
    process(i_clk)
        variable dx, dy     : integer;
        variable dist2      : integer;
        variable rad2       : integer := LED_RADIUS * LED_RADIUS;
        
        variable center_x   : integer;
        variable led_idx    : integer; -- 0 to 6
        variable is_led_on  : boolean;
        variable hit_circle : boolean;
        variable current_bit: std_logic;
    begin
        if rising_edge(i_clk) then
            if i_rst = '1' then
                o_red   <= (others => '0');
                o_green <= (others => '0');
                o_blue  <= (others => '0');
            elsif pix_ce = '1' then
                -- �w�]�I���� (�`�Ŧ�)
                o_red   <= "0000";
                o_green <= "0000";
                o_blue  <= "0010"; 
    
                if (h_count < H_RES) and (v_count < V_RES) then
                    hit_circle := false;
                    is_led_on  := false;
                    
                    -- �u�ơG���ˬd Y �b�O�_�b��νd�򤺡A��֭p��q
                    if abs(v_count - LED_Y) <= LED_RADIUS then
                        
                        -- �ˬd 7 �� LED ����m
                        -- �ڭ̰��] LED �q����k ���� led_status(6) �� led_status(0)
                        for k in 0 to 6 loop
                            center_x := LED_START_X + k * LED_GAP;
                            
                            -- �ˬd X �b�d�� (BBox check)
                            if abs(h_count - center_x) <= LED_RADIUS then
                                dx := h_count - center_x;
                                dy := v_count - LED_Y;
                                dist2 := dx*dx + dy*dy;
                                
                                if dist2 <= rad2 then
                                    hit_circle := true;
                                    
                                    -- ���� logic vector: �ù�����(k=0)���� Bit 6
                                    current_bit := led_status(6 - k);  -- �ھ� led_status �P�_�O�_��ܸ����y
                                    
                                    if current_bit = '1' then
                                        is_led_on := true;
                                    else
                                        is_led_on := false;
                                    end if;
                                    
                                    -- �ھ� led_status �]�w�C��
                                    if is_led_on then
                                        -- �ھ� led_status ��ܤ��P�C��
                                        case k is
                                            when 0 =>
                                                -- �C��]�w 1 (�Ҧp����)
                                                o_red   <= "1111";
                                                o_green <= "0000";
                                                o_blue  <= "0000";  -- Red
                                            when 1 =>
                                                -- �C��]�w 2 (�Ҧp���)
                                                o_red   <= "0000";
                                                o_green <= "1111";
                                                o_blue  <= "0000";  -- Green
                                            when 2 =>
                                                -- �C��]�w 3 (�Ҧp�Ŧ�)
                                                o_red   <= "0000";
                                                o_green <= "0000";
                                                o_blue  <= "1111";  -- Blue
                                            when 3 =>
                                                -- �C��]�w 4 (�Ҧp����)
                                                o_red   <= "1111";
                                                o_green <= "1111";
                                                o_blue  <= "0000";  -- Yellow
                                            when 4 =>
                                                -- �C��]�w 5 (�Ҧp����)
                                                o_red   <= "1111";
                                                o_green <= "0000";
                                                o_blue  <= "1111";  -- Purple
                                            when 5 =>
                                                -- �C��]�w 6 (�Ҧp�C��)
                                                o_red   <= "0000";
                                                o_green <= "1111";
                                                o_blue  <= "1111";  -- Cyan
                                            when 6 =>
                                                -- �C��]�w 7 (�Ҧp�զ�)
                                                o_red   <= "1111";
                                                o_green <= "1111";
                                                o_blue  <= "1111";  -- White
                                            when others =>
                                                -- ��L�C�� (�¦������)
                                                o_red   <= "0000";
                                                o_green <= "0000";
                                                o_blue  <= "0000";  -- Black or Off
                                        end case;
                                    else
                                        -- �p�G���� LED �S���Q�}�ҡA�h��ܭI���C��
                                        o_red   <= "0010";
                                        o_green <= "0010";
                                        o_blue  <= "0010";  -- Background (Blue)
                                    end if;
                                    
                                    -- ���@�Ӷ�N�����~���ˬd��L���F (�]���ꤣ���|)
                                    exit; 
                                end if;
                            end if;
                        end loop;
                        
                    end if; -- Y check
                else
                    -- Blanking Interval (�µe��)
                    o_red   <= (others => '0');
                    o_green <= (others => '0');
                    o_blue  <= (others => '0');
                end if;
            end if;
        end if;
    end process;
end rtl;
